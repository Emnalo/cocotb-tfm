module pic_rom (
    input [8:0] addr,
    output reg [11:0] data
);

    always @(*) begin
        case (addr)
            9'd0  : data = 12'b110000001001;
            9'd1  : data = 12'b000000101000;
            9'd2  : data = 12'b110000001000;
            9'd3  : data = 12'b000000101001;
            9'd4  : data = 12'b110000000111;
            9'd5  : data = 12'b000000101010;
            9'd6  : data = 12'b110000000110;
            9'd7  : data = 12'b000000101011;
            9'd8  : data = 12'b110000000101;
            9'd9  : data = 12'b000000101100;
            9'd10 : data = 12'b110000000100;
            9'd11 : data = 12'b000000101101;
            9'd12 : data = 12'b110000000011;
            9'd13 : data = 12'b000000101110;
            9'd14 : data = 12'b110000000010;
            9'd15 : data = 12'b000000101111;
            9'd16 : data = 12'b110000000001;
            9'd17 : data = 12'b000000110000;
            9'd18 : data = 12'b110000000000;
            9'd19 : data = 12'b000000110001;
            9'd20 : data = 12'b110000001000;
            9'd21 : data = 12'b000000100100;
            9'd22 : data = 12'b110000001001;
            9'd23 : data = 12'b000000110011;
            9'd24 : data = 12'b000111100100;
            9'd25 : data = 12'b001000000000;
            9'd26 : data = 12'b000000110010;
            9'd27 : data = 12'b000011100100;
            9'd28 : data = 12'b001000010010;
            9'd29 : data = 12'b000010000000;
            9'd30 : data = 12'b011101000011;
            9'd31 : data = 12'b101000100101;
            9'd32 : data = 12'b001000010010;
            9'd33 : data = 12'b000110100000;
            9'd34 : data = 12'b000110000000;
            9'd35 : data = 12'b000110100000;
            9'd36 : data = 12'b000000110010;
            9'd37 : data = 12'b110000001000;
            9'd38 : data = 12'b000110000100;
            9'd39 : data = 12'b011100000011;
            9'd40 : data = 12'b101000011011;
            9'd41 : data = 12'b110000001000;
            9'd42 : data = 12'b000111010011;
            9'd43 : data = 12'b000000100100;
            9'd44 : data = 12'b001000010010;
            9'd45 : data = 12'b000000100000;
            9'd46 : data = 12'b000011100100;
            9'd47 : data = 12'b001011110011;
            9'd48 : data = 12'b101000011001;
            9'd49 : data = 12'b000000000000;
            default: data = 12'b000000000000;
        endcase
    end

endmodule

