`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.08.2024 20:11:02
// Design Name: 
// Module Name: pic_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module pic_rom(
    input [8:0] Addr,
    output reg [11:0] Data
    );
    
    always @(Addr) begin
        case (Addr)
            0 : Data <= 12'b110000001001;
            1 : Data <= 12'b000000101000;
            2 : Data <= 12'b110000001000;
            3 : Data <= 12'b000000101001;
            4 : Data <= 12'b110000000111;
            5 : Data <= 12'b000000101010;
            6 : Data <= 12'b110000000110;
            7 : Data <= 12'b000000101011;
            8 : Data <= 12'b110000000101;
            9 : Data <= 12'b000000101100;
            10 : Data <= 12'b110000000100;
            11 : Data <= 12'b000000101101;
            12 : Data <= 12'b110000000011;
            13 : Data <= 12'b000000101110;
            14 : Data <= 12'b110000000010;
            15 : Data <= 12'b000000101111;
            16 : Data <= 12'b110000000001;
            17 : Data <= 12'b000000110000;
            18 : Data <= 12'b110000000000;
            19 : Data <= 12'b000000110001;
            20 : Data <= 12'b110000001000;
            21 : Data <= 12'b000000100100;
            22 : Data <= 12'b110000001001;
            23 : Data <= 12'b000000110011;
            24 : Data <= 12'b000111100100;
            25 : Data <= 12'b001000000000;
            26 : Data <= 12'b000000110010;
            27 : Data <= 12'b000011100100;
            28 : Data <= 12'b001000010010;
            29 : Data <= 12'b000010000000;
            30 : Data <= 12'b011101000011;
            31 : Data <= 12'b101000100101;
            32 : Data <= 12'b001000010010;
            33 : Data <= 12'b000110100000;
            34 : Data <= 12'b000110000000;
            35 : Data <= 12'b000110100000;
            36 : Data <= 12'b000000110010;
            37 : Data <= 12'b110000001000;
            38 : Data <= 12'b000110000100;
            39 : Data <= 12'b011100000011;
            40 : Data <= 12'b101000011011;
            41 : Data <= 12'b110000001000;
            42 : Data <= 12'b000111010011;
            43 : Data <= 12'b000000100100;
            44 : Data <= 12'b001000010010;
            45 : Data <= 12'b000000100000;
            46 : Data <= 12'b000011100100;
            47 : Data <= 12'b001011110011;
            48 : Data <= 12'b101000011001;
            default : Data <= 12'b000000000000;
        endcase
    end
    
endmodule
