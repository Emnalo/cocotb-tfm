library IEEE;
use IEEE.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.std_logic_arith.all;


entity ROM IS
  PORT (
    clk : IN STD_LOGIC;
    reset : IN STD_LOGIC;
    addr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    dout : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
        attribute bram_map: string;                     ---statement of the blockram
        attribute bram_map of ROM: entity is "yes";    
      
        attribute cascade_height : integer;
        attribute cascade_height of ROM: entity is 0;        
END ROM;





architecture Behavioral of ROM is

   type   memory is array (4095 downto 0) of std_logic_vector(7 downto 0);

    
    signal mem: memory := (
        0 => "00000010",
        1 => "00001010",
        2 => "11000110",
        3 => "00000000",
        4 => "00000000",
        5 => "00000000",
        6 => "00000000",
        7 => "00000000",
        8 => "00000000",
        9 => "00000000",
        10 => "00000000",
        11 => "00000000",
        12 => "00000000",
        13 => "00000000",
        14 => "00000000",
        15 => "00000000",
        16 => "00000000",
        17 => "00000000",
        18 => "00000000",
        19 => "00000000",
        20 => "00000000",
        21 => "00000000",
        22 => "00000000",
        23 => "00000000",
        24 => "00000000",
        25 => "00000000",
        26 => "00000000",
        27 => "00000000",
        28 => "00000000",
        29 => "00000000",
        30 => "00000000",
        31 => "00000000",
        32 => "00000000",
        33 => "00000000",
        34 => "00000000",
        35 => "00000000",
        36 => "00000000",
        37 => "00000000",
        38 => "00000000",
        39 => "00000000",
        40 => "00000000",
        41 => "00000000",
        42 => "00000000",
        43 => "00000000",
        44 => "00000000",
        45 => "00000000",
        46 => "00000000",
        47 => "00000000",
        48 => "00000000",
        49 => "00000000",
        50 => "00000000",
        51 => "00000000",
        52 => "00000000",
        53 => "00000000",
        54 => "00000000",
        55 => "00000000",
        56 => "00000000",
        57 => "00000000",
        58 => "00000000",
        59 => "00000000",
        60 => "00000000",
        61 => "00000000",
        62 => "00000000",
        63 => "00000000",
        64 => "00000000",
        65 => "00000000",
        66 => "00000000",
        67 => "00000000",
        68 => "00000000",
        69 => "00000000",
        70 => "00000000",
        71 => "00000000",
        72 => "00000000",
        73 => "00000000",
        74 => "00000000",
        75 => "00000000",
        76 => "00000000",
        77 => "00000000",
        78 => "00000000",
        79 => "00000000",
        80 => "00000000",
        81 => "00000000",
        82 => "00000000",
        83 => "00000000",
        84 => "00000000",
        85 => "00000000",
        86 => "00000000",
        87 => "00000000",
        88 => "00000000",
        89 => "00000000",
        90 => "00000000",
        91 => "00000000",
        92 => "00000000",
        93 => "00000000",
        94 => "00000000",
        95 => "00000000",
        96 => "00000000",
        97 => "00000000",
        98 => "00000000",
        99 => "00000000",
        100 => "00000000",
        101 => "00000000",
        102 => "00000000",
        103 => "00000000",
        104 => "00000000",
        105 => "00000000",
        106 => "00000000",
        107 => "00000000",
        108 => "00000000",
        109 => "00000000",
        110 => "00000000",
        111 => "00000000",
        112 => "00000000",
        113 => "00000000",
        114 => "00000000",
        115 => "00000000",
        116 => "00000000",
        117 => "00000000",
        118 => "00000000",
        119 => "00000000",
        120 => "00000000",
        121 => "00000000",
        122 => "00000000",
        123 => "00000000",
        124 => "00000000",
        125 => "00000000",
        126 => "00000000",
        127 => "00000000",
        128 => "00000000",
        129 => "00000000",
        130 => "00000000",
        131 => "00000000",
        132 => "00000000",
        133 => "00000000",
        134 => "00000000",
        135 => "00000000",
        136 => "00000000",
        137 => "00000000",
        138 => "00000000",
        139 => "00000000",
        140 => "00000000",
        141 => "00000000",
        142 => "00000000",
        143 => "00000000",
        144 => "00000000",
        145 => "00000000",
        146 => "00000000",
        147 => "00000000",
        148 => "00000000",
        149 => "00000000",
        150 => "00000000",
        151 => "00000000",
        152 => "00000000",
        153 => "00000000",
        154 => "00000000",
        155 => "00000000",
        156 => "00000000",
        157 => "00000000",
        158 => "00000000",
        159 => "00000000",
        160 => "00000000",
        161 => "00000000",
        162 => "00000000",
        163 => "00000000",
        164 => "00000000",
        165 => "00000000",
        166 => "00000000",
        167 => "00000000",
        168 => "00000000",
        169 => "00000000",
        170 => "00000000",
        171 => "00000000",
        172 => "00000000",
        173 => "00000000",
        174 => "00000000",
        175 => "00000000",
        176 => "00000000",
        177 => "00000000",
        178 => "00000000",
        179 => "00000000",
        180 => "00000000",
        181 => "00000000",
        182 => "00000000",
        183 => "00000000",
        184 => "00000000",
        185 => "00000000",
        186 => "00000000",
        187 => "00000000",
        188 => "00000000",
        189 => "00000000",
        190 => "00000000",
        191 => "00000000",
        192 => "00000000",
        193 => "00000000",
        194 => "00000000",
        195 => "00000000",
        196 => "00000000",
        197 => "00000000",
        198 => "00000000",
        199 => "00000000",
        200 => "00000000",
        201 => "00000000",
        202 => "00000000",
        203 => "00000000",
        204 => "00000000",
        205 => "00000000",
        206 => "00000000",
        207 => "00000000",
        208 => "00000000",
        209 => "00000000",
        210 => "00000000",
        211 => "00000000",
        212 => "00000000",
        213 => "00000000",
        214 => "00000000",
        215 => "00000000",
        216 => "00000000",
        217 => "00000000",
        218 => "00000000",
        219 => "00000000",
        220 => "00000000",
        221 => "00000000",
        222 => "00000000",
        223 => "00000000",
        224 => "00000000",
        225 => "00000000",
        226 => "00000000",
        227 => "00000000",
        228 => "00000000",
        229 => "00000000",
        230 => "00000000",
        231 => "00000000",
        232 => "00000000",
        233 => "00000000",
        234 => "00000000",
        235 => "00000000",
        236 => "00000000",
        237 => "00000000",
        238 => "00000000",
        239 => "00000000",
        240 => "00000000",
        241 => "00000000",
        242 => "00000000",
        243 => "00000000",
        244 => "00000000",
        245 => "00000000",
        246 => "00000000",
        247 => "00000000",
        248 => "00000000",
        249 => "00000000",
        250 => "00000000",
        251 => "00000000",
        252 => "00000000",
        253 => "00000000",
        254 => "00000000",
        255 => "00000000",
        256 => "00000000",
        257 => "00000000",
        258 => "00000000",
        259 => "00000000",
        260 => "00000000",
        261 => "00000000",
        262 => "00000000",
        263 => "00000000",
        264 => "00000000",
        265 => "00000000",
        266 => "00000000",
        267 => "00000000",
        268 => "00000000",
        269 => "00000000",
        270 => "00000000",
        271 => "00000000",
        272 => "00000000",
        273 => "00000000",
        274 => "00000000",
        275 => "00000000",
        276 => "00000000",
        277 => "00000000",
        278 => "00000000",
        279 => "00000000",
        280 => "00000000",
        281 => "00000000",
        282 => "00000000",
        283 => "00000000",
        284 => "00000000",
        285 => "00000000",
        286 => "00000000",
        287 => "00000000",
        288 => "00000000",
        289 => "00000000",
        290 => "00000000",
        291 => "00000000",
        292 => "00000000",
        293 => "00000000",
        294 => "00000000",
        295 => "00000000",
        296 => "00000000",
        297 => "00000000",
        298 => "00000000",
        299 => "00000000",
        300 => "00000000",
        301 => "00000000",
        302 => "00000000",
        303 => "00000000",
        304 => "00000000",
        305 => "00000000",
        306 => "00000000",
        307 => "00000000",
        308 => "00000000",
        309 => "00000000",
        310 => "00000000",
        311 => "00000000",
        312 => "00000000",
        313 => "00000000",
        314 => "00000000",
        315 => "00000000",
        316 => "00000000",
        317 => "00000000",
        318 => "00000000",
        319 => "00000000",
        320 => "00000000",
        321 => "00000000",
        322 => "00000000",
        323 => "00000000",
        324 => "00000000",
        325 => "00000000",
        326 => "00000000",
        327 => "00000000",
        328 => "00000000",
        329 => "00000000",
        330 => "00000000",
        331 => "00000000",
        332 => "00000000",
        333 => "00000000",
        334 => "00000000",
        335 => "00000000",
        336 => "00000000",
        337 => "00000000",
        338 => "00000000",
        339 => "00000000",
        340 => "00000000",
        341 => "00000000",
        342 => "00000000",
        343 => "00000000",
        344 => "00000000",
        345 => "00000000",
        346 => "00000000",
        347 => "00000000",
        348 => "00000000",
        349 => "00000000",
        350 => "00000000",
        351 => "00000000",
        352 => "00000000",
        353 => "00000000",
        354 => "00000000",
        355 => "00000000",
        356 => "00000000",
        357 => "00000000",
        358 => "00000000",
        359 => "00000000",
        360 => "00000000",
        361 => "00000000",
        362 => "00000000",
        363 => "00000000",
        364 => "00000000",
        365 => "00000000",
        366 => "00000000",
        367 => "00000000",
        368 => "00000000",
        369 => "00000000",
        370 => "00000000",
        371 => "00000000",
        372 => "00000000",
        373 => "00000000",
        374 => "00000000",
        375 => "00000000",
        376 => "00000000",
        377 => "00000000",
        378 => "00000000",
        379 => "00000000",
        380 => "00000000",
        381 => "00000000",
        382 => "00000000",
        383 => "00000000",
        384 => "00000000",
        385 => "00000000",
        386 => "00000000",
        387 => "00000000",
        388 => "00000000",
        389 => "00000000",
        390 => "00000000",
        391 => "00000000",
        392 => "00000000",
        393 => "00000000",
        394 => "00000000",
        395 => "00000000",
        396 => "00000000",
        397 => "00000000",
        398 => "00000000",
        399 => "00000000",
        400 => "00000000",
        401 => "00000000",
        402 => "00000000",
        403 => "00000000",
        404 => "00000000",
        405 => "00000000",
        406 => "00000000",
        407 => "00000000",
        408 => "00000000",
        409 => "00000000",
        410 => "00000000",
        411 => "00000000",
        412 => "00000000",
        413 => "00000000",
        414 => "00000000",
        415 => "00000000",
        416 => "00000000",
        417 => "00000000",
        418 => "00000000",
        419 => "00000000",
        420 => "00000000",
        421 => "00000000",
        422 => "00000000",
        423 => "00000000",
        424 => "00000000",
        425 => "00000000",
        426 => "00000000",
        427 => "00000000",
        428 => "00000000",
        429 => "00000000",
        430 => "00000000",
        431 => "00000000",
        432 => "00000000",
        433 => "00000000",
        434 => "00000000",
        435 => "00000000",
        436 => "00000000",
        437 => "00000000",
        438 => "00000000",
        439 => "00000000",
        440 => "00000000",
        441 => "00000000",
        442 => "00000000",
        443 => "00000000",
        444 => "00000000",
        445 => "00000000",
        446 => "00000000",
        447 => "00000000",
        448 => "00000000",
        449 => "00000000",
        450 => "00000000",
        451 => "00000000",
        452 => "00000000",
        453 => "00000000",
        454 => "00000000",
        455 => "00000000",
        456 => "00000000",
        457 => "00000000",
        458 => "00000000",
        459 => "00000000",
        460 => "00000000",
        461 => "00000000",
        462 => "00000000",
        463 => "00000000",
        464 => "00000000",
        465 => "00000000",
        466 => "00000000",
        467 => "00000000",
        468 => "00000000",
        469 => "00000000",
        470 => "00000000",
        471 => "00000000",
        472 => "00000000",
        473 => "00000000",
        474 => "00000000",
        475 => "00000000",
        476 => "00000000",
        477 => "00000000",
        478 => "00000000",
        479 => "00000000",
        480 => "00000000",
        481 => "00000000",
        482 => "00000000",
        483 => "00000000",
        484 => "00000000",
        485 => "00000000",
        486 => "00000000",
        487 => "00000000",
        488 => "00000000",
        489 => "00000000",
        490 => "00000000",
        491 => "00000000",
        492 => "00000000",
        493 => "00000000",
        494 => "00000000",
        495 => "00000000",
        496 => "00000000",
        497 => "00000000",
        498 => "00000000",
        499 => "00000000",
        500 => "00000000",
        501 => "00000000",
        502 => "00000000",
        503 => "00000000",
        504 => "00000000",
        505 => "00000000",
        506 => "00000000",
        507 => "00000000",
        508 => "00000000",
        509 => "00000000",
        510 => "00000000",
        511 => "00000000",
        512 => "00000000",
        513 => "00000000",
        514 => "00000000",
        515 => "00000000",
        516 => "00000000",
        517 => "00000000",
        518 => "00000000",
        519 => "00000000",
        520 => "00000000",
        521 => "00000000",
        522 => "00000000",
        523 => "00000000",
        524 => "00000000",
        525 => "00000000",
        526 => "00000000",
        527 => "00000000",
        528 => "00000000",
        529 => "00000000",
        530 => "00000000",
        531 => "00000000",
        532 => "00000000",
        533 => "00000000",
        534 => "00000000",
        535 => "00000000",
        536 => "00000000",
        537 => "00000000",
        538 => "00000000",
        539 => "00000000",
        540 => "00000000",
        541 => "00000000",
        542 => "00000000",
        543 => "00000000",
        544 => "00000000",
        545 => "00000000",
        546 => "00000000",
        547 => "00000000",
        548 => "00000000",
        549 => "00000000",
        550 => "00000000",
        551 => "00000000",
        552 => "00000000",
        553 => "00000000",
        554 => "00000000",
        555 => "00000000",
        556 => "00000000",
        557 => "00000000",
        558 => "00000000",
        559 => "00000000",
        560 => "00000000",
        561 => "00000000",
        562 => "00000000",
        563 => "00000000",
        564 => "00000000",
        565 => "00000000",
        566 => "00000000",
        567 => "00000000",
        568 => "00000000",
        569 => "00000000",
        570 => "00000000",
        571 => "00000000",
        572 => "00000000",
        573 => "00000000",
        574 => "00000000",
        575 => "00000000",
        576 => "00000000",
        577 => "00000000",
        578 => "00000000",
        579 => "00000000",
        580 => "00000000",
        581 => "00000000",
        582 => "00000000",
        583 => "00000000",
        584 => "00000000",
        585 => "00000000",
        586 => "00000000",
        587 => "00000000",
        588 => "00000000",
        589 => "00000000",
        590 => "00000000",
        591 => "00000000",
        592 => "00000000",
        593 => "00000000",
        594 => "00000000",
        595 => "00000000",
        596 => "00000000",
        597 => "00000000",
        598 => "00000000",
        599 => "00000000",
        600 => "00000000",
        601 => "00000000",
        602 => "00000000",
        603 => "00000000",
        604 => "00000000",
        605 => "00000000",
        606 => "00000000",
        607 => "00000000",
        608 => "00000000",
        609 => "00000000",
        610 => "00000000",
        611 => "00000000",
        612 => "00000000",
        613 => "00000000",
        614 => "00000000",
        615 => "00000000",
        616 => "00000000",
        617 => "00000000",
        618 => "00000000",
        619 => "00000000",
        620 => "00000000",
        621 => "00000000",
        622 => "00000000",
        623 => "00000000",
        624 => "00000000",
        625 => "00000000",
        626 => "00000000",
        627 => "00000000",
        628 => "00000000",
        629 => "00000000",
        630 => "00000000",
        631 => "00000000",
        632 => "00000000",
        633 => "00000000",
        634 => "00000000",
        635 => "00000000",
        636 => "00000000",
        637 => "00000000",
        638 => "00000000",
        639 => "00000000",
        640 => "00000000",
        641 => "00000000",
        642 => "00000000",
        643 => "00000000",
        644 => "00000000",
        645 => "00000000",
        646 => "00000000",
        647 => "00000000",
        648 => "00000000",
        649 => "00000000",
        650 => "00000000",
        651 => "00000000",
        652 => "00000000",
        653 => "00000000",
        654 => "00000000",
        655 => "00000000",
        656 => "00000000",
        657 => "00000000",
        658 => "00000000",
        659 => "00000000",
        660 => "00000000",
        661 => "00000000",
        662 => "00000000",
        663 => "00000000",
        664 => "00000000",
        665 => "00000000",
        666 => "00000000",
        667 => "00000000",
        668 => "00000000",
        669 => "00000000",
        670 => "00000000",
        671 => "00000000",
        672 => "00000000",
        673 => "00000000",
        674 => "00000000",
        675 => "00000000",
        676 => "00000000",
        677 => "00000000",
        678 => "00000000",
        679 => "00000000",
        680 => "00000000",
        681 => "00000000",
        682 => "00000000",
        683 => "00000000",
        684 => "00000000",
        685 => "00000000",
        686 => "00000000",
        687 => "00000000",
        688 => "00000000",
        689 => "00000000",
        690 => "00000000",
        691 => "00000000",
        692 => "00000000",
        693 => "00000000",
        694 => "00000000",
        695 => "00000000",
        696 => "00000000",
        697 => "00000000",
        698 => "00000000",
        699 => "00000000",
        700 => "00000000",
        701 => "00000000",
        702 => "00000000",
        703 => "00000000",
        704 => "00000000",
        705 => "00000000",
        706 => "00000000",
        707 => "00000000",
        708 => "00000000",
        709 => "00000000",
        710 => "00000000",
        711 => "00000000",
        712 => "00000000",
        713 => "00000000",
        714 => "00000000",
        715 => "00000000",
        716 => "00000000",
        717 => "00000000",
        718 => "00000000",
        719 => "00000000",
        720 => "00000000",
        721 => "00000000",
        722 => "00000000",
        723 => "00000000",
        724 => "00000000",
        725 => "00000000",
        726 => "00000000",
        727 => "00000000",
        728 => "00000000",
        729 => "00000000",
        730 => "00000000",
        731 => "00000000",
        732 => "00000000",
        733 => "00000000",
        734 => "00000000",
        735 => "00000000",
        736 => "00000000",
        737 => "00000000",
        738 => "00000000",
        739 => "00000000",
        740 => "00000000",
        741 => "00000000",
        742 => "00000000",
        743 => "00000000",
        744 => "00000000",
        745 => "00000000",
        746 => "00000000",
        747 => "00000000",
        748 => "00000000",
        749 => "00000000",
        750 => "00000000",
        751 => "00000000",
        752 => "00000000",
        753 => "00000000",
        754 => "00000000",
        755 => "00000000",
        756 => "00000000",
        757 => "00000000",
        758 => "00000000",
        759 => "00000000",
        760 => "00000000",
        761 => "00000000",
        762 => "00000000",
        763 => "00000000",
        764 => "00000000",
        765 => "00000000",
        766 => "00000000",
        767 => "00000000",
        768 => "00000000",
        769 => "00000000",
        770 => "00000000",
        771 => "00000000",
        772 => "00000000",
        773 => "00000000",
        774 => "00000000",
        775 => "00000000",
        776 => "00000000",
        777 => "00000000",
        778 => "00000000",
        779 => "00000000",
        780 => "00000000",
        781 => "00000000",
        782 => "00000000",
        783 => "00000000",
        784 => "00000000",
        785 => "00000000",
        786 => "00000000",
        787 => "00000000",
        788 => "00000000",
        789 => "00000000",
        790 => "00000000",
        791 => "00000000",
        792 => "00000000",
        793 => "00000000",
        794 => "00000000",
        795 => "00000000",
        796 => "00000000",
        797 => "00000000",
        798 => "00000000",
        799 => "00000000",
        800 => "00000000",
        801 => "00000000",
        802 => "00000000",
        803 => "00000000",
        804 => "00000000",
        805 => "00000000",
        806 => "00000000",
        807 => "00000000",
        808 => "00000000",
        809 => "00000000",
        810 => "00000000",
        811 => "00000000",
        812 => "00000000",
        813 => "00000000",
        814 => "00000000",
        815 => "00000000",
        816 => "00000000",
        817 => "00000000",
        818 => "00000000",
        819 => "00000000",
        820 => "00000000",
        821 => "00000000",
        822 => "00000000",
        823 => "00000000",
        824 => "00000000",
        825 => "00000000",
        826 => "00000000",
        827 => "00000000",
        828 => "00000000",
        829 => "00000000",
        830 => "00000000",
        831 => "00000000",
        832 => "00000000",
        833 => "00000000",
        834 => "00000000",
        835 => "00000000",
        836 => "00000000",
        837 => "00000000",
        838 => "00000000",
        839 => "00000000",
        840 => "00000000",
        841 => "00000000",
        842 => "00000000",
        843 => "00000000",
        844 => "00000000",
        845 => "00000000",
        846 => "00000000",
        847 => "00000000",
        848 => "00000000",
        849 => "00000000",
        850 => "00000000",
        851 => "00000000",
        852 => "00000000",
        853 => "00000000",
        854 => "00000000",
        855 => "00000000",
        856 => "00000000",
        857 => "00000000",
        858 => "00000000",
        859 => "00000000",
        860 => "00000000",
        861 => "00000000",
        862 => "00000000",
        863 => "00000000",
        864 => "00000000",
        865 => "00000000",
        866 => "00000000",
        867 => "00000000",
        868 => "00000000",
        869 => "00000000",
        870 => "00000000",
        871 => "00000000",
        872 => "00000000",
        873 => "00000000",
        874 => "00000000",
        875 => "00000000",
        876 => "00000000",
        877 => "00000000",
        878 => "00000000",
        879 => "00000000",
        880 => "00000000",
        881 => "00000000",
        882 => "00000000",
        883 => "00000000",
        884 => "00000000",
        885 => "00000000",
        886 => "00000000",
        887 => "00000000",
        888 => "00000000",
        889 => "00000000",
        890 => "00000000",
        891 => "00000000",
        892 => "00000000",
        893 => "00000000",
        894 => "00000000",
        895 => "00000000",
        896 => "00000000",
        897 => "00000000",
        898 => "00000000",
        899 => "00000000",
        900 => "00000000",
        901 => "00000000",
        902 => "00000000",
        903 => "00000000",
        904 => "00000000",
        905 => "00000000",
        906 => "00000000",
        907 => "00000000",
        908 => "00000000",
        909 => "00000000",
        910 => "00000000",
        911 => "00000000",
        912 => "00000000",
        913 => "00000000",
        914 => "00000000",
        915 => "00000000",
        916 => "00000000",
        917 => "00000000",
        918 => "00000000",
        919 => "00000000",
        920 => "00000000",
        921 => "00000000",
        922 => "00000000",
        923 => "00000000",
        924 => "00000000",
        925 => "00000000",
        926 => "00000000",
        927 => "00000000",
        928 => "00000000",
        929 => "00000000",
        930 => "00000000",
        931 => "00000000",
        932 => "00000000",
        933 => "00000000",
        934 => "00000000",
        935 => "00000000",
        936 => "00000000",
        937 => "00000000",
        938 => "00000000",
        939 => "00000000",
        940 => "00000000",
        941 => "00000000",
        942 => "00000000",
        943 => "00000000",
        944 => "00000000",
        945 => "00000000",
        946 => "00000000",
        947 => "00000000",
        948 => "00000000",
        949 => "00000000",
        950 => "00000000",
        951 => "00000000",
        952 => "00000000",
        953 => "00000000",
        954 => "00000000",
        955 => "00000000",
        956 => "00000000",
        957 => "00000000",
        958 => "00000000",
        959 => "00000000",
        960 => "00000000",
        961 => "00000000",
        962 => "00000000",
        963 => "00000000",
        964 => "00000000",
        965 => "00000000",
        966 => "00000000",
        967 => "00000000",
        968 => "00000000",
        969 => "00000000",
        970 => "00000000",
        971 => "00000000",
        972 => "00000000",
        973 => "00000000",
        974 => "00000000",
        975 => "00000000",
        976 => "00000000",
        977 => "00000000",
        978 => "00000000",
        979 => "00000000",
        980 => "00000000",
        981 => "00000000",
        982 => "00000000",
        983 => "00000000",
        984 => "00000000",
        985 => "00000000",
        986 => "00000000",
        987 => "00000000",
        988 => "00000000",
        989 => "00000000",
        990 => "00000000",
        991 => "00000000",
        992 => "00000000",
        993 => "00000000",
        994 => "00000000",
        995 => "00000000",
        996 => "00000000",
        997 => "00000000",
        998 => "00000000",
        999 => "00000000",
        1000 => "00000000",
        1001 => "00000000",
        1002 => "00000000",
        1003 => "00000000",
        1004 => "00000000",
        1005 => "00000000",
        1006 => "00000000",
        1007 => "00000000",
        1008 => "00000000",
        1009 => "00000000",
        1010 => "00000000",
        1011 => "00000000",
        1012 => "00000000",
        1013 => "00000000",
        1014 => "00000000",
        1015 => "00000000",
        1016 => "00000000",
        1017 => "00000000",
        1018 => "00000000",
        1019 => "00000000",
        1020 => "00000000",
        1021 => "00000000",
        1022 => "00000000",
        1023 => "00000000",
        1024 => "00000000",
        1025 => "00000000",
        1026 => "00000000",
        1027 => "00000000",
        1028 => "00000000",
        1029 => "00000000",
        1030 => "00000000",
        1031 => "00000000",
        1032 => "00000000",
        1033 => "00000000",
        1034 => "00000000",
        1035 => "00000000",
        1036 => "00000000",
        1037 => "00000000",
        1038 => "00000000",
        1039 => "00000000",
        1040 => "00000000",
        1041 => "00000000",
        1042 => "00000000",
        1043 => "00000000",
        1044 => "00000000",
        1045 => "00000000",
        1046 => "00000000",
        1047 => "00000000",
        1048 => "00000000",
        1049 => "00000000",
        1050 => "00000000",
        1051 => "00000000",
        1052 => "00000000",
        1053 => "00000000",
        1054 => "00000000",
        1055 => "00000000",
        1056 => "00000000",
        1057 => "00000000",
        1058 => "00000000",
        1059 => "00000000",
        1060 => "00000000",
        1061 => "00000000",
        1062 => "00000000",
        1063 => "00000000",
        1064 => "00000000",
        1065 => "00000000",
        1066 => "00000000",
        1067 => "00000000",
        1068 => "00000000",
        1069 => "00000000",
        1070 => "00000000",
        1071 => "00000000",
        1072 => "00000000",
        1073 => "00000000",
        1074 => "00000000",
        1075 => "00000000",
        1076 => "00000000",
        1077 => "00000000",
        1078 => "00000000",
        1079 => "00000000",
        1080 => "00000000",
        1081 => "00000000",
        1082 => "00000000",
        1083 => "00000000",
        1084 => "00000000",
        1085 => "00000000",
        1086 => "00000000",
        1087 => "00000000",
        1088 => "00000000",
        1089 => "00000000",
        1090 => "00000000",
        1091 => "00000000",
        1092 => "00000000",
        1093 => "00000000",
        1094 => "00000000",
        1095 => "00000000",
        1096 => "00000000",
        1097 => "00000000",
        1098 => "00000000",
        1099 => "00000000",
        1100 => "00000000",
        1101 => "00000000",
        1102 => "00000000",
        1103 => "00000000",
        1104 => "00000000",
        1105 => "00000000",
        1106 => "00000000",
        1107 => "00000000",
        1108 => "00000000",
        1109 => "00000000",
        1110 => "00000000",
        1111 => "00000000",
        1112 => "00000000",
        1113 => "00000000",
        1114 => "00000000",
        1115 => "00000000",
        1116 => "00000000",
        1117 => "00000000",
        1118 => "00000000",
        1119 => "00000000",
        1120 => "00000000",
        1121 => "00000000",
        1122 => "00000000",
        1123 => "00000000",
        1124 => "00000000",
        1125 => "00000000",
        1126 => "00000000",
        1127 => "00000000",
        1128 => "00000000",
        1129 => "00000000",
        1130 => "00000000",
        1131 => "00000000",
        1132 => "00000000",
        1133 => "00000000",
        1134 => "00000000",
        1135 => "00000000",
        1136 => "00000000",
        1137 => "00000000",
        1138 => "00000000",
        1139 => "00000000",
        1140 => "00000000",
        1141 => "00000000",
        1142 => "00000000",
        1143 => "00000000",
        1144 => "00000000",
        1145 => "00000000",
        1146 => "00000000",
        1147 => "00000000",
        1148 => "00000000",
        1149 => "00000000",
        1150 => "00000000",
        1151 => "00000000",
        1152 => "00000000",
        1153 => "00000000",
        1154 => "00000000",
        1155 => "00000000",
        1156 => "00000000",
        1157 => "00000000",
        1158 => "00000000",
        1159 => "00000000",
        1160 => "00000000",
        1161 => "00000000",
        1162 => "00000000",
        1163 => "00000000",
        1164 => "00000000",
        1165 => "00000000",
        1166 => "00000000",
        1167 => "00000000",
        1168 => "00000000",
        1169 => "00000000",
        1170 => "00000000",
        1171 => "00000000",
        1172 => "00000000",
        1173 => "00000000",
        1174 => "00000000",
        1175 => "00000000",
        1176 => "00000000",
        1177 => "00000000",
        1178 => "00000000",
        1179 => "00000000",
        1180 => "00000000",
        1181 => "00000000",
        1182 => "00000000",
        1183 => "00000000",
        1184 => "00000000",
        1185 => "00000000",
        1186 => "00000000",
        1187 => "00000000",
        1188 => "00000000",
        1189 => "00000000",
        1190 => "00000000",
        1191 => "00000000",
        1192 => "00000000",
        1193 => "00000000",
        1194 => "00000000",
        1195 => "00000000",
        1196 => "00000000",
        1197 => "00000000",
        1198 => "00000000",
        1199 => "00000000",
        1200 => "00000000",
        1201 => "00000000",
        1202 => "00000000",
        1203 => "00000000",
        1204 => "00000000",
        1205 => "00000000",
        1206 => "00000000",
        1207 => "00000000",
        1208 => "00000000",
        1209 => "00000000",
        1210 => "00000000",
        1211 => "00000000",
        1212 => "00000000",
        1213 => "00000000",
        1214 => "00000000",
        1215 => "00000000",
        1216 => "00000000",
        1217 => "00000000",
        1218 => "00000000",
        1219 => "00000000",
        1220 => "00000000",
        1221 => "00000000",
        1222 => "00000000",
        1223 => "00000000",
        1224 => "00000000",
        1225 => "00000000",
        1226 => "00000000",
        1227 => "00000000",
        1228 => "00000000",
        1229 => "00000000",
        1230 => "00000000",
        1231 => "00000000",
        1232 => "00000000",
        1233 => "00000000",
        1234 => "00000000",
        1235 => "00000000",
        1236 => "00000000",
        1237 => "00000000",
        1238 => "00000000",
        1239 => "00000000",
        1240 => "00000000",
        1241 => "00000000",
        1242 => "00000000",
        1243 => "00000000",
        1244 => "00000000",
        1245 => "00000000",
        1246 => "00000000",
        1247 => "00000000",
        1248 => "00000000",
        1249 => "00000000",
        1250 => "00000000",
        1251 => "00000000",
        1252 => "00000000",
        1253 => "00000000",
        1254 => "00000000",
        1255 => "00000000",
        1256 => "00000000",
        1257 => "00000000",
        1258 => "00000000",
        1259 => "00000000",
        1260 => "00000000",
        1261 => "00000000",
        1262 => "00000000",
        1263 => "00000000",
        1264 => "00000000",
        1265 => "00000000",
        1266 => "00000000",
        1267 => "00000000",
        1268 => "00000000",
        1269 => "00000000",
        1270 => "00000000",
        1271 => "00000000",
        1272 => "00000000",
        1273 => "00000000",
        1274 => "00000000",
        1275 => "00000000",
        1276 => "00000000",
        1277 => "00000000",
        1278 => "00000000",
        1279 => "00000000",
        1280 => "00000000",
        1281 => "00000000",
        1282 => "00000000",
        1283 => "00000000",
        1284 => "00000000",
        1285 => "00000000",
        1286 => "00000000",
        1287 => "00000000",
        1288 => "00000000",
        1289 => "00000000",
        1290 => "00000000",
        1291 => "00000000",
        1292 => "00000000",
        1293 => "00000000",
        1294 => "00000000",
        1295 => "00000000",
        1296 => "00000000",
        1297 => "00000000",
        1298 => "00000000",
        1299 => "00000000",
        1300 => "00000000",
        1301 => "00000000",
        1302 => "00000000",
        1303 => "00000000",
        1304 => "00000000",
        1305 => "00000000",
        1306 => "00000000",
        1307 => "00000000",
        1308 => "00000000",
        1309 => "00000000",
        1310 => "00000000",
        1311 => "00000000",
        1312 => "00000000",
        1313 => "00000000",
        1314 => "00000000",
        1315 => "00000000",
        1316 => "00000000",
        1317 => "00000000",
        1318 => "00000000",
        1319 => "00000000",
        1320 => "00000000",
        1321 => "00000000",
        1322 => "00000000",
        1323 => "00000000",
        1324 => "00000000",
        1325 => "00000000",
        1326 => "00000000",
        1327 => "00000000",
        1328 => "00000000",
        1329 => "00000000",
        1330 => "00000000",
        1331 => "00000000",
        1332 => "00000000",
        1333 => "00000000",
        1334 => "00000000",
        1335 => "00000000",
        1336 => "00000000",
        1337 => "00000000",
        1338 => "00000000",
        1339 => "00000000",
        1340 => "00000000",
        1341 => "00000000",
        1342 => "00000000",
        1343 => "00000000",
        1344 => "00000000",
        1345 => "00000000",
        1346 => "00000000",
        1347 => "00000000",
        1348 => "00000000",
        1349 => "00000000",
        1350 => "00000000",
        1351 => "00000000",
        1352 => "00000000",
        1353 => "00000000",
        1354 => "00000000",
        1355 => "00000000",
        1356 => "00000000",
        1357 => "00000000",
        1358 => "00000000",
        1359 => "00000000",
        1360 => "00000000",
        1361 => "00000000",
        1362 => "00000000",
        1363 => "00000000",
        1364 => "00000000",
        1365 => "00000000",
        1366 => "00000000",
        1367 => "00000000",
        1368 => "00000000",
        1369 => "00000000",
        1370 => "00000000",
        1371 => "00000000",
        1372 => "00000000",
        1373 => "00000000",
        1374 => "00000000",
        1375 => "00000000",
        1376 => "00000000",
        1377 => "00000000",
        1378 => "00000000",
        1379 => "00000000",
        1380 => "00000000",
        1381 => "00000000",
        1382 => "00000000",
        1383 => "00000000",
        1384 => "00000000",
        1385 => "00000000",
        1386 => "00000000",
        1387 => "00000000",
        1388 => "00000000",
        1389 => "00000000",
        1390 => "00000000",
        1391 => "00000000",
        1392 => "00000000",
        1393 => "00000000",
        1394 => "00000000",
        1395 => "00000000",
        1396 => "00000000",
        1397 => "00000000",
        1398 => "00000000",
        1399 => "00000000",
        1400 => "00000000",
        1401 => "00000000",
        1402 => "00000000",
        1403 => "00000000",
        1404 => "00000000",
        1405 => "00000000",
        1406 => "00000000",
        1407 => "00000000",
        1408 => "00000000",
        1409 => "00000000",
        1410 => "00000000",
        1411 => "00000000",
        1412 => "00000000",
        1413 => "00000000",
        1414 => "00000000",
        1415 => "00000000",
        1416 => "00000000",
        1417 => "00000000",
        1418 => "00000000",
        1419 => "00000000",
        1420 => "00000000",
        1421 => "00000000",
        1422 => "00000000",
        1423 => "00000000",
        1424 => "00000000",
        1425 => "00000000",
        1426 => "00000000",
        1427 => "00000000",
        1428 => "00000000",
        1429 => "00000000",
        1430 => "00000000",
        1431 => "00000000",
        1432 => "00000000",
        1433 => "00000000",
        1434 => "00000000",
        1435 => "00000000",
        1436 => "00000000",
        1437 => "00000000",
        1438 => "00000000",
        1439 => "00000000",
        1440 => "00000000",
        1441 => "00000000",
        1442 => "00000000",
        1443 => "00000000",
        1444 => "00000000",
        1445 => "00000000",
        1446 => "00000000",
        1447 => "00000000",
        1448 => "00000000",
        1449 => "00000000",
        1450 => "00000000",
        1451 => "00000000",
        1452 => "00000000",
        1453 => "00000000",
        1454 => "00000000",
        1455 => "00000000",
        1456 => "00000000",
        1457 => "00000000",
        1458 => "00000000",
        1459 => "00000000",
        1460 => "00000000",
        1461 => "00000000",
        1462 => "00000000",
        1463 => "00000000",
        1464 => "00000000",
        1465 => "00000000",
        1466 => "00000000",
        1467 => "00000000",
        1468 => "00000000",
        1469 => "00000000",
        1470 => "00000000",
        1471 => "00000000",
        1472 => "00000000",
        1473 => "00000000",
        1474 => "00000000",
        1475 => "00000000",
        1476 => "00000000",
        1477 => "00000000",
        1478 => "00000000",
        1479 => "00000000",
        1480 => "00000000",
        1481 => "00000000",
        1482 => "00000000",
        1483 => "00000000",
        1484 => "00000000",
        1485 => "00000000",
        1486 => "00000000",
        1487 => "00000000",
        1488 => "00000000",
        1489 => "00000000",
        1490 => "00000000",
        1491 => "00000000",
        1492 => "00000000",
        1493 => "00000000",
        1494 => "00000000",
        1495 => "00000000",
        1496 => "00000000",
        1497 => "00000000",
        1498 => "00000000",
        1499 => "00000000",
        1500 => "00000000",
        1501 => "00000000",
        1502 => "00000000",
        1503 => "00000000",
        1504 => "00000000",
        1505 => "00000000",
        1506 => "00000000",
        1507 => "00000000",
        1508 => "00000000",
        1509 => "00000000",
        1510 => "00000000",
        1511 => "00000000",
        1512 => "00000000",
        1513 => "00000000",
        1514 => "00000000",
        1515 => "00000000",
        1516 => "00000000",
        1517 => "00000000",
        1518 => "00000000",
        1519 => "00000000",
        1520 => "00000000",
        1521 => "00000000",
        1522 => "00000000",
        1523 => "00000000",
        1524 => "00000000",
        1525 => "00000000",
        1526 => "00000000",
        1527 => "00000000",
        1528 => "00000000",
        1529 => "00000000",
        1530 => "00000000",
        1531 => "00000000",
        1532 => "00000000",
        1533 => "00000000",
        1534 => "00000000",
        1535 => "00000000",
        1536 => "00000000",
        1537 => "00000000",
        1538 => "00000000",
        1539 => "00000000",
        1540 => "00000000",
        1541 => "00000000",
        1542 => "00000000",
        1543 => "00000000",
        1544 => "00000000",
        1545 => "00000000",
        1546 => "00000000",
        1547 => "00000000",
        1548 => "00000000",
        1549 => "00000000",
        1550 => "00000000",
        1551 => "00000000",
        1552 => "00000000",
        1553 => "00000000",
        1554 => "00000000",
        1555 => "00000000",
        1556 => "00000000",
        1557 => "00000000",
        1558 => "00000000",
        1559 => "00000000",
        1560 => "00000000",
        1561 => "00000000",
        1562 => "00000000",
        1563 => "00000000",
        1564 => "00000000",
        1565 => "00000000",
        1566 => "00000000",
        1567 => "00000000",
        1568 => "00000000",
        1569 => "00000000",
        1570 => "00000000",
        1571 => "00000000",
        1572 => "00000000",
        1573 => "00000000",
        1574 => "00000000",
        1575 => "00000000",
        1576 => "00000000",
        1577 => "00000000",
        1578 => "00000000",
        1579 => "00000000",
        1580 => "00000000",
        1581 => "00000000",
        1582 => "00000000",
        1583 => "00000000",
        1584 => "00000000",
        1585 => "00000000",
        1586 => "00000000",
        1587 => "00000000",
        1588 => "00000000",
        1589 => "00000000",
        1590 => "00000000",
        1591 => "00000000",
        1592 => "00000000",
        1593 => "00000000",
        1594 => "00000000",
        1595 => "00000000",
        1596 => "00000000",
        1597 => "00000000",
        1598 => "00000000",
        1599 => "00000000",
        1600 => "00000000",
        1601 => "00000000",
        1602 => "00000000",
        1603 => "00000000",
        1604 => "00000000",
        1605 => "00000000",
        1606 => "00000000",
        1607 => "00000000",
        1608 => "00000000",
        1609 => "00000000",
        1610 => "00000000",
        1611 => "00000000",
        1612 => "00000000",
        1613 => "00000000",
        1614 => "00000000",
        1615 => "00000000",
        1616 => "00000000",
        1617 => "00000000",
        1618 => "00000000",
        1619 => "00000000",
        1620 => "00000000",
        1621 => "00000000",
        1622 => "00000000",
        1623 => "00000000",
        1624 => "00000000",
        1625 => "00000000",
        1626 => "00000000",
        1627 => "00000000",
        1628 => "00000000",
        1629 => "00000000",
        1630 => "00000000",
        1631 => "00000000",
        1632 => "00000000",
        1633 => "00000000",
        1634 => "00000000",
        1635 => "00000000",
        1636 => "00000000",
        1637 => "00000000",
        1638 => "00000000",
        1639 => "00000000",
        1640 => "00000000",
        1641 => "00000000",
        1642 => "00000000",
        1643 => "00000000",
        1644 => "00000000",
        1645 => "00000000",
        1646 => "00000000",
        1647 => "00000000",
        1648 => "00000000",
        1649 => "00000000",
        1650 => "00000000",
        1651 => "00000000",
        1652 => "00000000",
        1653 => "00000000",
        1654 => "00000000",
        1655 => "00000000",
        1656 => "00000000",
        1657 => "00000000",
        1658 => "00000000",
        1659 => "00000000",
        1660 => "00000000",
        1661 => "00000000",
        1662 => "00000000",
        1663 => "00000000",
        1664 => "00000000",
        1665 => "00000000",
        1666 => "00000000",
        1667 => "00000000",
        1668 => "00000000",
        1669 => "00000000",
        1670 => "00000000",
        1671 => "00000000",
        1672 => "00000000",
        1673 => "00000000",
        1674 => "00000000",
        1675 => "00000000",
        1676 => "00000000",
        1677 => "00000000",
        1678 => "00000000",
        1679 => "00000000",
        1680 => "00000000",
        1681 => "00000000",
        1682 => "00000000",
        1683 => "00000000",
        1684 => "00000000",
        1685 => "00000000",
        1686 => "00000000",
        1687 => "00000000",
        1688 => "00000000",
        1689 => "00000000",
        1690 => "00000000",
        1691 => "00000000",
        1692 => "00000000",
        1693 => "00000000",
        1694 => "00000000",
        1695 => "00000000",
        1696 => "00000000",
        1697 => "00000000",
        1698 => "00000000",
        1699 => "00000000",
        1700 => "00000000",
        1701 => "00000000",
        1702 => "00000000",
        1703 => "00000000",
        1704 => "00000000",
        1705 => "00000000",
        1706 => "00000000",
        1707 => "00000000",
        1708 => "00000000",
        1709 => "00000000",
        1710 => "00000000",
        1711 => "00000000",
        1712 => "00000000",
        1713 => "00000000",
        1714 => "00000000",
        1715 => "00000000",
        1716 => "00000000",
        1717 => "00000000",
        1718 => "00000000",
        1719 => "00000000",
        1720 => "00000000",
        1721 => "00000000",
        1722 => "00000000",
        1723 => "00000000",
        1724 => "00000000",
        1725 => "00000000",
        1726 => "00000000",
        1727 => "00000000",
        1728 => "00000000",
        1729 => "00000000",
        1730 => "00000000",
        1731 => "00000000",
        1732 => "00000000",
        1733 => "00000000",
        1734 => "00000000",
        1735 => "00000000",
        1736 => "00000000",
        1737 => "00000000",
        1738 => "00000000",
        1739 => "00000000",
        1740 => "00000000",
        1741 => "00000000",
        1742 => "00000000",
        1743 => "00000000",
        1744 => "00000000",
        1745 => "00000000",
        1746 => "00000000",
        1747 => "00000000",
        1748 => "00000000",
        1749 => "00000000",
        1750 => "00000000",
        1751 => "00000000",
        1752 => "00000000",
        1753 => "00000000",
        1754 => "00000000",
        1755 => "00000000",
        1756 => "00000000",
        1757 => "00000000",
        1758 => "00000000",
        1759 => "00000000",
        1760 => "00000000",
        1761 => "00000000",
        1762 => "00000000",
        1763 => "00000000",
        1764 => "00000000",
        1765 => "00000000",
        1766 => "00000000",
        1767 => "00000000",
        1768 => "00000000",
        1769 => "00000000",
        1770 => "00000000",
        1771 => "00000000",
        1772 => "00000000",
        1773 => "00000000",
        1774 => "00000000",
        1775 => "00000000",
        1776 => "00000000",
        1777 => "00000000",
        1778 => "00000000",
        1779 => "00000000",
        1780 => "00000000",
        1781 => "00000000",
        1782 => "00000000",
        1783 => "00000000",
        1784 => "00000000",
        1785 => "00000000",
        1786 => "00000000",
        1787 => "00000000",
        1788 => "00000000",
        1789 => "00000000",
        1790 => "00000000",
        1791 => "00000000",
        1792 => "00000000",
        1793 => "00000000",
        1794 => "00000000",
        1795 => "00000000",
        1796 => "00000000",
        1797 => "00000000",
        1798 => "00000000",
        1799 => "00000000",
        1800 => "00000000",
        1801 => "00000000",
        1802 => "00000000",
        1803 => "00000000",
        1804 => "00000000",
        1805 => "00000000",
        1806 => "00000000",
        1807 => "00000000",
        1808 => "00000000",
        1809 => "00000000",
        1810 => "00000000",
        1811 => "00000000",
        1812 => "00000000",
        1813 => "00000000",
        1814 => "00000000",
        1815 => "00000000",
        1816 => "00000000",
        1817 => "00000000",
        1818 => "00000000",
        1819 => "00000000",
        1820 => "00000000",
        1821 => "00000000",
        1822 => "00000000",
        1823 => "00000000",
        1824 => "00000000",
        1825 => "00000000",
        1826 => "00000000",
        1827 => "00000000",
        1828 => "00000000",
        1829 => "00000000",
        1830 => "00000000",
        1831 => "00000000",
        1832 => "00000000",
        1833 => "00000000",
        1834 => "00000000",
        1835 => "00000000",
        1836 => "00000000",
        1837 => "00000000",
        1838 => "00000000",
        1839 => "00000000",
        1840 => "00000000",
        1841 => "00000000",
        1842 => "00000000",
        1843 => "00000000",
        1844 => "00000000",
        1845 => "00000000",
        1846 => "00000000",
        1847 => "00000000",
        1848 => "00000000",
        1849 => "00000000",
        1850 => "00000000",
        1851 => "00000000",
        1852 => "00000000",
        1853 => "00000000",
        1854 => "00000000",
        1855 => "00000000",
        1856 => "00000000",
        1857 => "00000000",
        1858 => "00000000",
        1859 => "00000000",
        1860 => "00000000",
        1861 => "00000000",
        1862 => "00000000",
        1863 => "00000000",
        1864 => "00000000",
        1865 => "00000000",
        1866 => "00000000",
        1867 => "00000000",
        1868 => "00000000",
        1869 => "00000000",
        1870 => "00000000",
        1871 => "00000000",
        1872 => "00000000",
        1873 => "00000000",
        1874 => "00000000",
        1875 => "00000000",
        1876 => "00000000",
        1877 => "00000000",
        1878 => "00000000",
        1879 => "00000000",
        1880 => "00000000",
        1881 => "00000000",
        1882 => "00000000",
        1883 => "00000000",
        1884 => "00000000",
        1885 => "00000000",
        1886 => "00000000",
        1887 => "00000000",
        1888 => "00000000",
        1889 => "00000000",
        1890 => "00000000",
        1891 => "00000000",
        1892 => "00000000",
        1893 => "00000000",
        1894 => "00000000",
        1895 => "00000000",
        1896 => "00000000",
        1897 => "00000000",
        1898 => "00000000",
        1899 => "00000000",
        1900 => "00000000",
        1901 => "00000000",
        1902 => "00000000",
        1903 => "00000000",
        1904 => "00000000",
        1905 => "00000000",
        1906 => "00000000",
        1907 => "00000000",
        1908 => "00000000",
        1909 => "00000000",
        1910 => "00000000",
        1911 => "00000000",
        1912 => "00000000",
        1913 => "00000000",
        1914 => "00000000",
        1915 => "00000000",
        1916 => "00000000",
        1917 => "00000000",
        1918 => "00000000",
        1919 => "00000000",
        1920 => "00000000",
        1921 => "00000000",
        1922 => "00000000",
        1923 => "00000000",
        1924 => "00000000",
        1925 => "00000000",
        1926 => "00000000",
        1927 => "00000000",
        1928 => "00000000",
        1929 => "00000000",
        1930 => "00000000",
        1931 => "00000000",
        1932 => "00000000",
        1933 => "00000000",
        1934 => "00000000",
        1935 => "00000000",
        1936 => "00000000",
        1937 => "00000000",
        1938 => "00000000",
        1939 => "00000000",
        1940 => "00000000",
        1941 => "00000000",
        1942 => "00000000",
        1943 => "00000000",
        1944 => "00000000",
        1945 => "00000000",
        1946 => "00000000",
        1947 => "00000000",
        1948 => "00000000",
        1949 => "00000000",
        1950 => "00000000",
        1951 => "00000000",
        1952 => "00000000",
        1953 => "00000000",
        1954 => "00000000",
        1955 => "00000000",
        1956 => "00000000",
        1957 => "00000000",
        1958 => "00000000",
        1959 => "00000000",
        1960 => "00000000",
        1961 => "00000000",
        1962 => "00000000",
        1963 => "00000000",
        1964 => "00000000",
        1965 => "00000000",
        1966 => "00000000",
        1967 => "00000000",
        1968 => "00000000",
        1969 => "00000000",
        1970 => "00000000",
        1971 => "00000000",
        1972 => "00000000",
        1973 => "00000000",
        1974 => "00000000",
        1975 => "00000000",
        1976 => "00000000",
        1977 => "00000000",
        1978 => "00000000",
        1979 => "00000000",
        1980 => "00000000",
        1981 => "00000000",
        1982 => "00000000",
        1983 => "00000000",
        1984 => "00000000",
        1985 => "00000000",
        1986 => "00000000",
        1987 => "00000000",
        1988 => "00000000",
        1989 => "00000000",
        1990 => "00000000",
        1991 => "00000000",
        1992 => "00000000",
        1993 => "00000000",
        1994 => "00000000",
        1995 => "00000000",
        1996 => "00000000",
        1997 => "00000000",
        1998 => "00000000",
        1999 => "00000000",
        2000 => "00000000",
        2001 => "00000000",
        2002 => "00000000",
        2003 => "00000000",
        2004 => "00000000",
        2005 => "00000000",
        2006 => "00000000",
        2007 => "00000000",
        2008 => "00000000",
        2009 => "00000000",
        2010 => "00000000",
        2011 => "00000000",
        2012 => "00000000",
        2013 => "00000000",
        2014 => "00000000",
        2015 => "00000000",
        2016 => "00000000",
        2017 => "00000000",
        2018 => "00000000",
        2019 => "00000000",
        2020 => "00000000",
        2021 => "00000000",
        2022 => "00000000",
        2023 => "00000000",
        2024 => "00000000",
        2025 => "00000000",
        2026 => "00000000",
        2027 => "00000000",
        2028 => "00000000",
        2029 => "00000000",
        2030 => "00000000",
        2031 => "00000000",
        2032 => "00000000",
        2033 => "00000000",
        2034 => "00000000",
        2035 => "00000000",
        2036 => "00000000",
        2037 => "00000000",
        2038 => "00000000",
        2039 => "00000000",
        2040 => "00000000",
        2041 => "00000000",
        2042 => "00000000",
        2043 => "00000000",
        2044 => "00000000",
        2045 => "00000000",
        2046 => "00000000",
        2047 => "00000000",
        2048 => "11100100",
        2049 => "11110101",
        2050 => "00001110",
        2051 => "11110101",
        2052 => "00001111",
        2053 => "01110101",
        2054 => "00010000",
        2055 => "00000001",
        2056 => "01110101",
        2057 => "00010001",
        2058 => "00000000",
        2059 => "01110101",
        2060 => "00010010",
        2061 => "00000000",
        2062 => "11110101",
        2063 => "00001000",
        2064 => "11110101",
        2065 => "00001001",
        2066 => "11100100",
        2067 => "11110101",
        2068 => "00001010",
        2069 => "11110101",
        2070 => "00001011",
        2071 => "11100101",
        2072 => "00001011",
        2073 => "00100101",
        2074 => "11100000",
        2075 => "11111111",
        2076 => "11100101",
        2077 => "00001010",
        2078 => "00110011",
        2079 => "11111110",
        2080 => "10010000",
        2081 => "00000000",
        2082 => "00000000",
        2083 => "01110101",
        2084 => "11110000",
        2085 => "00001010",
        2086 => "11100101",
        2087 => "00001001",
        2088 => "00010010",
        2089 => "00001010",
        2090 => "00011101",
        2091 => "11100101",
        2092 => "00001000",
        2093 => "01110101",
        2094 => "11110000",
        2095 => "00001010",
        2096 => "10100100",
        2097 => "00100101",
        2098 => "10000011",
        2099 => "11110101",
        2100 => "10000011",
        2101 => "11100101",
        2102 => "10000010",
        2103 => "00101111",
        2104 => "11110101",
        2105 => "10000010",
        2106 => "11100101",
        2107 => "10000011",
        2108 => "00111110",
        2109 => "11110101",
        2110 => "10000011",
        2111 => "11100100",
        2112 => "11110000",
        2113 => "10100011",
        2114 => "11110000",
        2115 => "11110101",
        2116 => "00001100",
        2117 => "11110101",
        2118 => "00001101",
        2119 => "11100101",
        2120 => "00001101",
        2121 => "00100101",
        2122 => "11100000",
        2123 => "11111101",
        2124 => "11100101",
        2125 => "00001100",
        2126 => "00110011",
        2127 => "11111100",
        2128 => "11100101",
        2129 => "00001001",
        2130 => "10101110",
        2131 => "00001000",
        2132 => "01111000",
        2133 => "00000011",
        2134 => "11000011",
        2135 => "00110011",
        2136 => "11001110",
        2137 => "00110011",
        2138 => "11001110",
        2139 => "11011000",
        2140 => "11111001",
        2141 => "00100100",
        2142 => "01111110",
        2143 => "11110101",
        2144 => "10000010",
        2145 => "01110100",
        2146 => "00001010",
        2147 => "00111110",
        2148 => "11110101",
        2149 => "10000011",
        2150 => "11100101",
        2151 => "10000010",
        2152 => "00101101",
        2153 => "11110101",
        2154 => "10000010",
        2155 => "11100101",
        2156 => "10000011",
        2157 => "00111100",
        2158 => "11110101",
        2159 => "10000011",
        2160 => "11100100",
        2161 => "10010011",
        2162 => "11111010",
        2163 => "01110100",
        2164 => "00000001",
        2165 => "10010011",
        2166 => "11111011",
        2167 => "11100101",
        2168 => "00001011",
        2169 => "00100101",
        2170 => "11100000",
        2171 => "11111111",
        2172 => "11100101",
        2173 => "00001010",
        2174 => "00110011",
        2175 => "11111110",
        2176 => "10010000",
        2177 => "00001010",
        2178 => "10011110",
        2179 => "01110101",
        2180 => "11110000",
        2181 => "00001010",
        2182 => "11100101",
        2183 => "00001101",
        2184 => "00010010",
        2185 => "00001010",
        2186 => "00011101",
        2187 => "11100101",
        2188 => "00001100",
        2189 => "01110101",
        2190 => "11110000",
        2191 => "00001010",
        2192 => "10100100",
        2193 => "00100101",
        2194 => "10000011",
        2195 => "11110101",
        2196 => "10000011",
        2197 => "11100101",
        2198 => "10000010",
        2199 => "00101111",
        2200 => "11110101",
        2201 => "10000010",
        2202 => "11100101",
        2203 => "10000011",
        2204 => "00111110",
        2205 => "11110101",
        2206 => "10000011",
        2207 => "11100100",
        2208 => "10010011",
        2209 => "11111100",
        2210 => "01110100",
        2211 => "00000001",
        2212 => "10010011",
        2213 => "11111101",
        2214 => "10101111",
        2215 => "00000011",
        2216 => "10101110",
        2217 => "00000010",
        2218 => "00010010",
        2219 => "00001001",
        2220 => "10000111",
        2221 => "10101100",
        2222 => "00000110",
        2223 => "10101101",
        2224 => "00000111",
        2225 => "11100101",
        2226 => "00001011",
        2227 => "00100101",
        2228 => "11100000",
        2229 => "11111111",
        2230 => "11100101",
        2231 => "00001010",
        2232 => "00110011",
        2233 => "11111110",
        2234 => "10010000",
        2235 => "00000000",
        2236 => "00000000",
        2237 => "01110101",
        2238 => "11110000",
        2239 => "00001010",
        2240 => "11100101",
        2241 => "00001001",
        2242 => "00010010",
        2243 => "00001010",
        2244 => "00011101",
        2245 => "11100101",
        2246 => "00001000",
        2247 => "01110101",
        2248 => "11110000",
        2249 => "00001010",
        2250 => "10100100",
        2251 => "00100101",
        2252 => "10000011",
        2253 => "11110101",
        2254 => "10000011",
        2255 => "11100101",
        2256 => "10000010",
        2257 => "00101111",
        2258 => "11110101",
        2259 => "10000010",
        2260 => "11100101",
        2261 => "10000011",
        2262 => "00111110",
        2263 => "11110101",
        2264 => "10000011",
        2265 => "11101100",
        2266 => "10001101",
        2267 => "11110000",
        2268 => "00010010",
        2269 => "00001001",
        2270 => "11001111",
        2271 => "00000101",
        2272 => "00001101",
        2273 => "11100101",
        2274 => "00001101",
        2275 => "01110000",
        2276 => "00000010",
        2277 => "00000101",
        2278 => "00001100",
        2279 => "01100100",
        2280 => "00000100",
        2281 => "01000101",
        2282 => "00001100",
        2283 => "01100000",
        2284 => "00000011",
        2285 => "00000010",
        2286 => "00001000",
        2287 => "01000111",
        2288 => "00000101",
        2289 => "00001011",
        2290 => "11100101",
        2291 => "00001011",
        2292 => "01110000",
        2293 => "00000010",
        2294 => "00000101",
        2295 => "00001010",
        2296 => "01100100",
        2297 => "00000101",
        2298 => "01000101",
        2299 => "00001010",
        2300 => "01100000",
        2301 => "00000011",
        2302 => "00000010",
        2303 => "00001000",
        2304 => "00010111",
        2305 => "00000101",
        2306 => "00001001",
        2307 => "11100101",
        2308 => "00001001",
        2309 => "01110000",
        2310 => "00000010",
        2311 => "00000101",
        2312 => "00001000",
        2313 => "01100100",
        2314 => "00000100",
        2315 => "01000101",
        2316 => "00001000",
        2317 => "01100000",
        2318 => "00000011",
        2319 => "00000010",
        2320 => "00001000",
        2321 => "00010010",
        2322 => "11100100",
        2323 => "11110101",
        2324 => "00001010",
        2325 => "11110101",
        2326 => "00001011",
        2327 => "11100101",
        2328 => "00001011",
        2329 => "00100101",
        2330 => "11100000",
        2331 => "11111011",
        2332 => "11100101",
        2333 => "00001010",
        2334 => "00110011",
        2335 => "11111010",
        2336 => "01110100",
        2337 => "00000000",
        2338 => "00101011",
        2339 => "11110101",
        2340 => "10000010",
        2341 => "01110100",
        2342 => "00000000",
        2343 => "00111010",
        2344 => "11110101",
        2345 => "10000011",
        2346 => "11100000",
        2347 => "11111110",
        2348 => "10100011",
        2349 => "11100000",
        2350 => "11111111",
        2351 => "10101101",
        2352 => "10000000",
        2353 => "11101101",
        2354 => "00100100",
        2355 => "00000001",
        2356 => "11111101",
        2357 => "11100100",
        2358 => "00110011",
        2359 => "11111100",
        2360 => "00010010",
        2361 => "00001001",
        2362 => "10011001",
        2363 => "10101101",
        2364 => "10000000",
        2365 => "11101111",
        2366 => "01001101",
        2367 => "11111111",
        2368 => "01110100",
        2369 => "00000000",
        2370 => "00101011",
        2371 => "11110101",
        2372 => "10000010",
        2373 => "01110100",
        2374 => "00000000",
        2375 => "00111010",
        2376 => "11110101",
        2377 => "10000011",
        2378 => "11101110",
        2379 => "11110000",
        2380 => "10100011",
        2381 => "11101111",
        2382 => "11110000",
        2383 => "00000101",
        2384 => "00001011",
        2385 => "11100101",
        2386 => "00001011",
        2387 => "01110000",
        2388 => "00000010",
        2389 => "00000101",
        2390 => "00001010",
        2391 => "01100100",
        2392 => "00000101",
        2393 => "01000101",
        2394 => "00001010",
        2395 => "01110000",
        2396 => "10111010",
        2397 => "11100101",
        2398 => "00001111",
        2399 => "00100101",
        2400 => "11100000",
        2401 => "11111111",
        2402 => "11100101",
        2403 => "00001110",
        2404 => "00110011",
        2405 => "10101011",
        2406 => "00010000",
        2407 => "10101010",
        2408 => "00010001",
        2409 => "10101001",
        2410 => "00010010",
        2411 => "10001111",
        2412 => "10000010",
        2413 => "11110101",
        2414 => "10000011",
        2415 => "00010010",
        2416 => "00001001",
        2417 => "11100101",
        2418 => "11110101",
        2419 => "00010100",
        2420 => "10000101",
        2421 => "11110000",
        2422 => "00010011",
        2423 => "11110101",
        2424 => "10010000",
        2425 => "11100101",
        2426 => "00010011",
        2427 => "11111111",
        2428 => "10001111",
        2429 => "10100000",
        2430 => "10101111",
        2431 => "10110000",
        2432 => "01110101",
        2433 => "00001110",
        2434 => "00000000",
        2435 => "10001111",
        2436 => "00001111",
        2437 => "10000000",
        2438 => "11010110",
        2439 => "11101111",
        2440 => "10001101",
        2441 => "11110000",
        2442 => "10100100",
        2443 => "10101000",
        2444 => "11110000",
        2445 => "11001111",
        2446 => "10001100",
        2447 => "11110000",
        2448 => "10100100",
        2449 => "00101000",
        2450 => "11001110",
        2451 => "10001101",
        2452 => "11110000",
        2453 => "10100100",
        2454 => "00101110",
        2455 => "11111110",
        2456 => "00100010",
        2457 => "11000010",
        2458 => "11010101",
        2459 => "11101100",
        2460 => "00110000",
        2461 => "11100111",
        2462 => "00001001",
        2463 => "10110010",
        2464 => "11010101",
        2465 => "11100100",
        2466 => "11000011",
        2467 => "10011101",
        2468 => "11111101",
        2469 => "11100100",
        2470 => "10011100",
        2471 => "11111100",
        2472 => "11101110",
        2473 => "00110000",
        2474 => "11100111",
        2475 => "00010101",
        2476 => "10110010",
        2477 => "11010101",
        2478 => "11100100",
        2479 => "11000011",
        2480 => "10011111",
        2481 => "11111111",
        2482 => "11100100",
        2483 => "10011110",
        2484 => "11111110",
        2485 => "00010010",
        2486 => "00001010",
        2487 => "00101001",
        2488 => "11000011",
        2489 => "11100100",
        2490 => "10011101",
        2491 => "11111101",
        2492 => "11100100",
        2493 => "10011100",
        2494 => "11111100",
        2495 => "10000000",
        2496 => "00000011",
        2497 => "00010010",
        2498 => "00001010",
        2499 => "00101001",
        2500 => "00110000",
        2501 => "11010101",
        2502 => "00000111",
        2503 => "11000011",
        2504 => "11100100",
        2505 => "10011111",
        2506 => "11111111",
        2507 => "11100100",
        2508 => "10011110",
        2509 => "11111110",
        2510 => "00100010",
        2511 => "11000101",
        2512 => "11110000",
        2513 => "11111000",
        2514 => "10100011",
        2515 => "11100000",
        2516 => "00101000",
        2517 => "11110000",
        2518 => "11000101",
        2519 => "11110000",
        2520 => "11111000",
        2521 => "11100101",
        2522 => "10000010",
        2523 => "00010101",
        2524 => "10000010",
        2525 => "01110000",
        2526 => "00000010",
        2527 => "00010101",
        2528 => "10000011",
        2529 => "11100000",
        2530 => "00111000",
        2531 => "11110000",
        2532 => "00100010",
        2533 => "10111011",
        2534 => "00000001",
        2535 => "00010000",
        2536 => "11100101",
        2537 => "10000010",
        2538 => "00101001",
        2539 => "11110101",
        2540 => "10000010",
        2541 => "11100101",
        2542 => "10000011",
        2543 => "00111010",
        2544 => "11110101",
        2545 => "10000011",
        2546 => "11100000",
        2547 => "11110101",
        2548 => "11110000",
        2549 => "10100011",
        2550 => "11100000",
        2551 => "00100010",
        2552 => "01010000",
        2553 => "00001001",
        2554 => "11101001",
        2555 => "00100101",
        2556 => "10000010",
        2557 => "11111000",
        2558 => "10000110",
        2559 => "11110000",
        2560 => "00001000",
        2561 => "11100110",
        2562 => "00100010",
        2563 => "10111011",
        2564 => "11111110",
        2565 => "00001010",
        2566 => "11101001",
        2567 => "00100101",
        2568 => "10000010",
        2569 => "11111000",
        2570 => "11100010",
        2571 => "11110101",
        2572 => "11110000",
        2573 => "00001000",
        2574 => "11100010",
        2575 => "00100010",
        2576 => "11100101",
        2577 => "10000011",
        2578 => "00101010",
        2579 => "11110101",
        2580 => "10000011",
        2581 => "11101001",
        2582 => "10010011",
        2583 => "11110101",
        2584 => "11110000",
        2585 => "10100011",
        2586 => "11101001",
        2587 => "10010011",
        2588 => "00100010",
        2589 => "10100100",
        2590 => "00100101",
        2591 => "10000010",
        2592 => "11110101",
        2593 => "10000010",
        2594 => "11100101",
        2595 => "11110000",
        2596 => "00110101",
        2597 => "10000011",
        2598 => "11110101",
        2599 => "10000011",
        2600 => "00100010",
        2601 => "10111100",
        2602 => "00000000",
        2603 => "00001011",
        2604 => "10111110",
        2605 => "00000000",
        2606 => "00101001",
        2607 => "11101111",
        2608 => "10001101",
        2609 => "11110000",
        2610 => "10000100",
        2611 => "11111111",
        2612 => "10101101",
        2613 => "11110000",
        2614 => "00100010",
        2615 => "11100100",
        2616 => "11001100",
        2617 => "11111000",
        2618 => "01110101",
        2619 => "11110000",
        2620 => "00001000",
        2621 => "11101111",
        2622 => "00101111",
        2623 => "11111111",
        2624 => "11101110",
        2625 => "00110011",
        2626 => "11111110",
        2627 => "11101100",
        2628 => "00110011",
        2629 => "11111100",
        2630 => "11101110",
        2631 => "10011101",
        2632 => "11101100",
        2633 => "10011000",
        2634 => "01000000",
        2635 => "00000101",
        2636 => "11111100",
        2637 => "11101110",
        2638 => "10011101",
        2639 => "11111110",
        2640 => "00001111",
        2641 => "11010101",
        2642 => "11110000",
        2643 => "11101001",
        2644 => "11100100",
        2645 => "11001110",
        2646 => "11111101",
        2647 => "00100010",
        2648 => "11101101",
        2649 => "11111000",
        2650 => "11110101",
        2651 => "11110000",
        2652 => "11101110",
        2653 => "10000100",
        2654 => "00100000",
        2655 => "11010010",
        2656 => "00011100",
        2657 => "11111110",
        2658 => "10101101",
        2659 => "11110000",
        2660 => "01110101",
        2661 => "11110000",
        2662 => "00001000",
        2663 => "11101111",
        2664 => "00101111",
        2665 => "11111111",
        2666 => "11101101",
        2667 => "00110011",
        2668 => "11111101",
        2669 => "01000000",
        2670 => "00000111",
        2671 => "10011000",
        2672 => "01010000",
        2673 => "00000110",
        2674 => "11010101",
        2675 => "11110000",
        2676 => "11110010",
        2677 => "00100010",
        2678 => "11000011",
        2679 => "10011000",
        2680 => "11111101",
        2681 => "00001111",
        2682 => "11010101",
        2683 => "11110000",
        2684 => "11101010",
        2685 => "00100010",
        2686 => "00010011",
        2687 => "00111111",
        2688 => "11011110",
        2689 => "01011100",
        2690 => "01101110",
        2691 => "10000010",
        2692 => "11110000",
        2693 => "10001110",
        2694 => "11000100",
        2695 => "10000010",
        2696 => "00000000",
        2697 => "00000111",
        2698 => "11010010",
        2699 => "01110101",
        2700 => "01001100",
        2701 => "10010000",
        2702 => "11101001",
        2703 => "01010101",
        2704 => "11111111",
        2705 => "11110010",
        2706 => "00100101",
        2707 => "00111101",
        2708 => "11111100",
        2709 => "01101101",
        2710 => "01001110",
        2711 => "10010011",
        2712 => "00001110",
        2713 => "11000111",
        2714 => "11100010",
        2715 => "11010011",
        2716 => "00000011",
        2717 => "11111111",
        2718 => "11010011",
        2719 => "00100100",
        2720 => "00001111",
        2721 => "10100000",
        2722 => "00000000",
        2723 => "01001111",
        2724 => "00011100",
        2725 => "10001111",
        2726 => "00000001",
        2727 => "00000000",
        2728 => "01001100",
        2729 => "10001110",
        2730 => "00000001",
        2731 => "11110111",
        2732 => "00000010",
        2733 => "10100010",
        2734 => "10000010",
        2735 => "00101110",
        2736 => "00001111",
        2737 => "10101010",
        2738 => "00100101",
        2739 => "01101100",
        2740 => "11111111",
        2741 => "10010101",
        2742 => "11111100",
        2743 => "11011000",
        2744 => "11101110",
        2745 => "10000101",
        2746 => "11111101",
        2747 => "01110000",
        2748 => "11111111",
        2749 => "11111111",
        2750 => "11111111",
        2751 => "11011001",
        2752 => "00000000",
        2753 => "10000000",
        2754 => "00000111",
        2755 => "00000001",
        2756 => "11111111",
        2757 => "00000001",
        2758 => "01111000",
        2759 => "01111111",
        2760 => "11100100",
        2761 => "11110110",
        2762 => "11011000",
        2763 => "11111101",
        2764 => "01110101",
        2765 => "10000001",
        2766 => "00010100",
        2767 => "00000010",
        2768 => "00001000",
        others => "00000000"    
    );
    

   
   
   attribute ram_style        : string;
   attribute ram_style of mem : signal is "block";  

   attribute cascade_height of mem: signal is 0;

   
   signal outreg : std_logic_vector(7 downto 0);

begin
       dout <= outreg  when reset='0'  else "00000000";

        process (clk)
            begin
              if (clk'event and clk='1') then
                if(addr(15 downto 12) = "0000") then 
                    outreg <= mem(conv_integer(unsigned(addr(11 downto 0)))); 
                else   
                    outreg <= "00000000";
                end if;
              end if;
        end process; 
  
end Behavioral;