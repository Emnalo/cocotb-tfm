`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.08.2024 20:11:02
// Design Name: 
// Module Name: pic_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module pic_rom(
    input [8:0] addr,
    output reg [11:0] data
    );
    
    always @(addr) begin
        case (addr)
            0 : data <= 12'b110000001001;
            1 : data <= 12'b000000101000;
            2 : data <= 12'b110000001000;
            3 : data <= 12'b000000101001;
            4 : data <= 12'b110000000111;
            5 : data <= 12'b000000101010;
            6 : data <= 12'b110000000110;
            7 : data <= 12'b000000101011;
            8 : data <= 12'b110000000101;
            9 : data <= 12'b000000101100;
            10 : data <= 12'b110000000100;
            11 : data <= 12'b000000101101;
            12 : data <= 12'b110000000011;
            13 : data <= 12'b000000101110;
            14 : data <= 12'b110000000010;
            15 : data <= 12'b000000101111;
            16 : data <= 12'b110000000001;
            17 : data <= 12'b000000110000;
            18 : data <= 12'b110000000000;
            19 : data <= 12'b000000110001;
            20 : data <= 12'b110000001000;
            21 : data <= 12'b000000100100;
            22 : data <= 12'b110000001001;
            23 : data <= 12'b000000110011;
            24 : data <= 12'b000111100100;
            25 : data <= 12'b001000000000;
            26 : data <= 12'b000000110010;
            27 : data <= 12'b000011100100;
            28 : data <= 12'b001000010010;
            29 : data <= 12'b000010000000;
            30 : data <= 12'b011101000011;
            31 : data <= 12'b101000100101;
            32 : data <= 12'b001000010010;
            33 : data <= 12'b000110100000;
            34 : data <= 12'b000110000000;
            35 : data <= 12'b000110100000;
            36 : data <= 12'b000000110010;
            37 : data <= 12'b110000001000;
            38 : data <= 12'b000110000100;
            39 : data <= 12'b011100000011;
            40 : data <= 12'b101000011011;
            41 : data <= 12'b110000001000;
            42 : data <= 12'b000111010011;
            43 : data <= 12'b000000100100;
            44 : data <= 12'b001000010010;
            45 : data <= 12'b000000100000;
            46 : data <= 12'b000011100100;
            47 : data <= 12'b001011110011;
            48 : data <= 12'b101000011001;
            default : data <= 12'b000000000000;
        endcase
    end
    
endmodule
